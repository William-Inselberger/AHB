module instructionmemory(
input [9:0]pc,
output reg [22:0]instruction
);


reg [22:0] memoria [0:1023];
integer i;
initial begin

	// WRITE_BURST(XXX)_SEL_ADDR(XX_XXXX_XXXX)_DATA(XXXX_XXXX)
	// write : 2 clk
	//read: 5 clk
	  
		memoria[0]=23'b0_000_0_00_0000_0000_0000_0000;  
    	memoria[1]=23'b1_000_0_00_0000_0001_0000_0001;  //1
		memoria[2]=23'b0_000_0_00_0000_0001_0000_0000; 
		memoria[3]=23'b1_000_0_00_0000_0010_0000_0010;	//2
		memoria[4]=23'b0_000_0_00_0000_0010_0000_0000;
		memoria[5]=23'b1_000_0_00_0000_0011_0000_0011;  //3
		memoria[6]=23'b0_000_0_00_0000_0011_0000_0000;
		memoria[7]=23'b1_000_0_00_0000_0100_0000_0100;  //4
		memoria[8]=23'b0_000_0_00_0000_0100_0000_0000;
		memoria[9]=23'b1_000_0_00_0000_0101_0000_0101;	//5
		memoria[10]=23'b0_000_0_00_0000_0101_0000_0000;
		memoria[11]=23'b1_000_0_00_0000_0110_0000_0110;	//6
		memoria[12]=23'b0_000_0_00_0000_0110_0000_0000;
		memoria[13]=23'b1_000_0_00_0000_0111_0000_0111; //7
		memoria[14]=23'b0_000_0_00_0000_0111_0000_0000;
		memoria[15]=23'b1_000_0_00_0000_1000_0000_1000; //8
		memoria[16]=23'b0_000_0_00_0000_1000_0000_0000;
		memoria[17]=23'b1_000_0_00_0000_1001_0000_1001; //9
		memoria[18]=23'b0_000_0_00_0000_1001_0000_0000;
		memoria[19]=23'b1_000_0_00_0000_1010_0000_1010;	//10
		memoria[20]=23'b0_000_0_00_0000_1010_0000_0000;
		memoria[21]=23'b1_000_0_00_0000_1011_0000_1011; //11
		memoria[22]=23'b0_000_0_00_0000_1011_0000_0000;
		
		memoria[23]=23'b0_000_1_00_0000_0000_0000_0000;  
    	memoria[24]=23'b1_000_1_00_0000_0001_0001_0001; //17
		memoria[25]=23'b0_000_1_00_0000_0001_0000_0000; 
		memoria[26]=23'b1_000_1_00_0000_0010_0001_0010; //18
		memoria[27]=23'b0_000_1_00_0000_0010_0000_0000;
		memoria[28]=23'b1_000_1_00_0000_0011_0001_0011; //19
		memoria[29]=23'b0_000_1_00_0000_0011_0000_0000;
		memoria[30]=23'b1_000_1_00_0000_0100_0001_0100; //20
		memoria[31]=23'b0_000_1_00_0000_0100_0000_0000;
		memoria[32]=23'b1_000_1_00_0000_0101_0001_0101; //21
		memoria[33]=23'b0_000_1_00_0000_0101_0000_0000;
		memoria[34]=23'b1_000_1_00_0000_0110_0001_0110; //22
		memoria[35]=23'b0_000_1_00_0000_0110_0000_0000;
		memoria[36]=23'b1_000_1_00_0000_0111_0001_0111; //23
		memoria[37]=23'b0_000_1_00_0000_0111_0000_0000;
		memoria[38]=23'b1_000_1_00_0000_1000_0001_1000; //24
		memoria[39]=23'b0_000_1_00_0000_1000_0000_0000;
		memoria[40]=23'b1_000_1_00_0000_1001_0001_1001; //25
		memoria[41]=23'b0_000_1_00_0000_1001_0000_0000;
		memoria[42]=23'b1_000_1_00_0000_1010_0001_1010; //26
		memoria[43]=23'b0_000_1_00_0000_1010_0000_0000;
		memoria[44]=23'b1_000_1_00_0000_1011_0001_1011; //27
		memoria[45]=23'b0_000_1_00_0000_1011_0000_0000;
	
end


always @(pc) begin

instruction = memoria[pc];

end







endmodule

